library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.DigEng.ALL; -- allows use of logarithms
-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity param_ALU_tb is
--  testbench empty entity
end param_ALU_tb;


architecture Behavioral of param_ALU_tb is
    constant data_size : NATURAL := 16;
    signal A : STD_LOGIC_VECTOR (data_size -1 downto 0);
    signal B : STD_LOGIC_VECTOR (data_size -1 downto 0);
    signal opcode : STD_LOGIC_VECTOR (3 downto 0);
    signal SH : UNSIGNED (log2(data_size)-1 downto 0); -- shift address
    signal Output : STD_LOGIC_VECTOR (data_size -1 downto 0); -- ALU output of [data_size] bits
    signal flags : STD_LOGIC_VECTOR(7 downto 0); -- flags encoded in fixed 8-bit bus
    
    type test_vector is record
        A_TV : STD_LOGIC_VECTOR (data_size-1 downto 0);
        B_TV : STD_LOGIC_VECTOR (data_size-1 downto 0);
        opcode_TV : STD_LOGIC_VECTOR (3 downto 0);   
        SH_TV :  UNSIGNED (log2(data_size)-1 downto 0);
        Output_TV : STD_LOGIC_VECTOR (data_size -1 downto 0);
        flags_TV : STD_LOGIC_VECTOR(7 downto 0);
    end record;
    
        
        
    type test_vector_array is array (NATURAL range <>) of test_vector;
            
    constant test_vectors : test_vector_array := (
        --Identity ALU_OUT <= A
        --[0, 32767, -32768, 1, -6550, -8876, 12079, -13440, 18614, 14010]
        (b"0000000000000000", b"0000000000000000", b"0000", b"0000", b"0000000000000000", b"01100001"),
        (b"0111111111111111", b"0000000000000000", b"0000", b"0000", b"0111111111111111", b"01010010"),
        (b"1000000000000000", b"0000000000000000", b"0000", b"0000", b"1000000000000000", b"00101010"),
        (b"0000000000000001", b"0000000000000000", b"0000", b"0000", b"0000000000000001", b"01010110"),
        (b"1110011001101010", b"0000000000000000", b"0000", b"0000", b"1110011001101010", b"00101010"),
        (b"1101110101010100", b"0000000000000000", b"0000", b"0000", b"1101110101010100", b"00101010"),
        (b"0010111100101111", b"0000000000000000", b"0000", b"0000", b"0010111100101111", b"01010010"),
        (b"1100101110000000", b"0000000000000000", b"0000", b"0000", b"1100101110000000", b"00101010"),
        (b"0100100010110110", b"0000000000000000", b"0000", b"0000", b"0100100010110110", b"01010010"),
        (b"0011011010111010", b"0000000000000000", b"0000", b"0000", b"0011011010111010", b"01010010"),
        --A&B
        --[0, 32767, -32768, 1, -12904, 27332, 1111, 15745, -31199, -4998, 1915, 15607, 14296, 27785, 5845]
        --[31300, 32183, -16853, -19143, -10608, 91, -23965, 10978, 23024, -25186, 15213, -2283, -12679, -5167, 10282]
        (b"0000000000000000", b"0111101001000100", b"0100", b"0000", b"0000000000000000", b"01100001"),
        (b"0111111111111111", b"0111110110110111", b"0100", b"0000", b"0111110110110111", b"01010010"),
        (b"1000000000000000", b"1011111000101011", b"0100", b"0000", b"1000000000000000", b"00101010"),
        (b"0000000000000001", b"1011010100111001", b"0100", b"0000", b"0000000000000001", b"01010110"),
        (b"1100110110011000", b"1101011010010000", b"0100", b"0000", b"1100010010010000", b"00101010"),
        (b"0110101011000100", b"0000000001011011", b"0100", b"0000", b"0000000001000000", b"01010010"),
        (b"0000010001010111", b"1010001001100011", b"0100", b"0000", b"0000000001000011", b"01010010"),
        (b"0011110110000001", b"0010101011100010", b"0100", b"0000", b"0010100010000000", b"01010010"),
        (b"1000011000100001", b"0101100111110000", b"0100", b"0000", b"0000000000100000", b"01010010"),
        (b"1110110001111010", b"1001110110011110", b"0100", b"0000", b"1000110000011010", b"00101010"),
        (b"0000011101111011", b"0011101101101101", b"0100", b"0000", b"0000001101101001", b"01010010"),
        (b"0011110011110111", b"1111011100010101", b"0100", b"0000", b"0011010000010101", b"01010010"),
        (b"0011011111011000", b"1100111001111001", b"0100", b"0000", b"0000011001011000", b"01010010"),
        (b"0110110010001001", b"1110101111010001", b"0100", b"0000", b"0110100010000001", b"01010010"),
        (b"0001011011010101", b"0010100000101010", b"0100", b"0000", b"0000000000000000", b"01100001"),
        --A | B
        --[0, 32767, -32768, 1, 26316, 28487, -857, -13317, -9269, 21998, -6751, 8094, -28005, -27492, -31845]
        --[32669, -9161, 26818, 17261, 9919, 27840, -5921, 15627, 16319, 22929, 17657, 7203, -23328, 5690, 10024]
        (b"0000000000000000", b"0111111110011101", b"0101", b"0000", b"0111111110011101", b"01010010"),
        (b"0111111111111111", b"1101110000110111", b"0101", b"0000", b"1111111111111111", b"00101010"),
        (b"1000000000000000", b"0110100011000010", b"0101", b"0000", b"1110100011000010", b"00101010"),
        (b"0000000000000001", b"0100001101101101", b"0101", b"0000", b"0100001101101101", b"01010010"),
        (b"0110011011001100", b"0010011010111111", b"0101", b"0000", b"0110011011111111", b"01010010"),
        (b"0110111101000111", b"0110110011000000", b"0101", b"0000", b"0110111111000111", b"01010010"),
        (b"1111110010100111", b"1110100011011111", b"0101", b"0000", b"1111110011111111", b"00101010"),
        (b"1100101111111011", b"0011110100001011", b"0101", b"0000", b"1111111111111011", b"00101010"),
        (b"1101101111001011", b"0011111110111111", b"0101", b"0000", b"1111111111111111", b"00101010"),
        (b"0101010111101110", b"0101100110010001", b"0101", b"0000", b"0101110111111111", b"01010010"),
        (b"1110010110100001", b"0100010011111001", b"0101", b"0000", b"1110010111111001", b"00101010"),
        (b"0001111110011110", b"0001110000100011", b"0101", b"0000", b"0001111110111111", b"01010010"),
        (b"1001001010011011", b"1010010011100000", b"0101", b"0000", b"1011011011111011", b"00101010"),
        (b"1001010010011100", b"0001011000111010", b"0101", b"0000", b"1001011010111110", b"00101010"),
        (b"1000001110011011", b"0010011100101000", b"0101", b"0000", b"1010011110111011", b"00101010"),
        --A XOR B 
        --[0, 32767, -32768, 1, 18164, 14065, -21984, -4590, 15337, -23716, -21644, 23269, -9070, 2620, -475]
        --[24459, 30605, 170, -3236, 31813, -23333, 18460, 30551, 19902, 22032, 32634, 2263, -8577, 394, 12874]
        (b"0000000000000000", b"0101111110001011", b"0110", b"0000", b"0101111110001011", b"01010010"),
        (b"0111111111111111", b"0111011110001101", b"0110", b"0000", b"0000100001110010", b"01010010"),
        (b"1000000000000000", b"0000000010101010", b"0110", b"0000", b"1000000010101010", b"00101010"),
        (b"0000000000000001", b"1111001101011100", b"0110", b"0000", b"1111001101011101", b"00101010"),
        (b"0100011011110100", b"0111110001000101", b"0110", b"0000", b"0011101010110001", b"01010010"),
        (b"0011011011110001", b"1010010011011011", b"0110", b"0000", b"1001001000101010", b"00101010"),
        (b"1010101000100000", b"0100100000011100", b"0110", b"0000", b"1110001000111100", b"00101010"),
        (b"1110111000010010", b"0111011101010111", b"0110", b"0000", b"1001100101000101", b"00101010"),
        (b"0011101111101001", b"0100110110111110", b"0110", b"0000", b"0111011001010111", b"01010010"),
        (b"1010001101011100", b"0101011000010000", b"0110", b"0000", b"1111010101001100", b"00101010"),
        (b"1010101101110100", b"0111111101111010", b"0110", b"0000", b"1101010000001110", b"00101010"),
        (b"0101101011100101", b"0000100011010111", b"0110", b"0000", b"0101001000110010", b"01010010"),
        (b"1101110010010010", b"1101111001111111", b"0110", b"0000", b"0000001011101101", b"01010010"),
        (b"0000101000111100", b"0000000110001010", b"0110", b"0000", b"0000101110110110", b"01010010"),
        (b"1111111000100101", b"0011001001001010", b"0110", b"0000", b"1100110001101111", b"00101010"),
        --NOT A
        --[0, 32767, -32768, 1, -5406, -30712, -22895, 32504, -27286, 15071, 14827, -1983, 412, 9756, -10817]
        --[0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0]
        (b"0000000000000000", b"0000000000000000", b"0111", b"0000", b"1111111111111111", b"00101010"),
        (b"0111111111111111", b"0000000000000000", b"0111", b"0000", b"1000000000000000", b"00101010"),
        (b"1000000000000000", b"0000000000000000", b"0111", b"0000", b"0111111111111111", b"01010010"),
        (b"0000000000000001", b"0000000000000000", b"0111", b"0000", b"1111111111111110", b"00101010"),
        (b"1110101011100010", b"0000000000000000", b"0111", b"0000", b"0001010100011101", b"01010010"),
        (b"1000100000001000", b"0000000000000000", b"0111", b"0000", b"0111011111110111", b"01010010"),
        (b"1010011010010001", b"0000000000000000", b"0111", b"0000", b"0101100101101110", b"01010010"),
        (b"0111111011111000", b"0000000000000000", b"0111", b"0000", b"1000000100000111", b"00101010"),
        (b"1001010101101010", b"0000000000000000", b"0111", b"0000", b"0110101010010101", b"01010010"),
        (b"0011101011011111", b"0000000000000000", b"0111", b"0000", b"1100010100100000", b"00101010"),
        (b"0011100111101011", b"0000000000000000", b"0111", b"0000", b"1100011000010100", b"00101010"),
        (b"1111100001000001", b"0000000000000000", b"0111", b"0000", b"0000011110111110", b"01010010"),
        (b"0000000110011100", b"0000000000000000", b"0111", b"0000", b"1111111001100011", b"00101010"),
        (b"0010011000011100", b"0000000000000000", b"0111", b"0000", b"1101100111100011", b"00101010"),
        (b"1101010110111111", b"0000000000000000", b"0111", b"0000", b"0010101001000000", b"01010010"),
        --A+1
        --[0, 32767, -32768, 1, 963, 2426, -7829, -1238, 23762, -13571, 26011, -15780, -18491, 16297, 28820]
        --[0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0]
        (b"0000000000000000", b"0000000000000000", b"1000", b"0000", b"0000000000000001", b"01010110"),
        (b"0111111111111111", b"0000000000000000", b"1000", b"0000", b"1000000000000000", b"11010010"),
        (b"1000000000000000", b"0000000000000000", b"1000", b"0000", b"1000000000000001", b"00101010"),
        (b"0000000000000001", b"0000000000000000", b"1000", b"0000", b"0000000000000010", b"01010010"),
        (b"0000001111000011", b"0000000000000000", b"1000", b"0000", b"0000001111000100", b"01010010"),
        (b"0000100101111010", b"0000000000000000", b"1000", b"0000", b"0000100101111011", b"01010010"),
        (b"1110000101101011", b"0000000000000000", b"1000", b"0000", b"1110000101101100", b"00101010"),
        (b"1111101100101010", b"0000000000000000", b"1000", b"0000", b"1111101100101011", b"00101010"),
        (b"0101110011010010", b"0000000000000000", b"1000", b"0000", b"0101110011010011", b"01010010"),
        (b"1100101011111101", b"0000000000000000", b"1000", b"0000", b"1100101011111110", b"00101010"),
        (b"0110010110011011", b"0000000000000000", b"1000", b"0000", b"0110010110011100", b"01010010"),
        (b"1100001001011100", b"0000000000000000", b"1000", b"0000", b"1100001001011101", b"00101010"),
        (b"1011011111000101", b"0000000000000000", b"1000", b"0000", b"1011011111000110", b"00101010"),
        (b"0011111110101001", b"0000000000000000", b"1000", b"0000", b"0011111110101010", b"01010010"),
        (b"0111000010010100", b"0000000000000000", b"1000", b"0000", b"0111000010010101", b"01010010"),
        --A-1
        --[0, 32767, -32768, 1, -11988, -22295, 22814, -18631, 29350, 15169, 3346, -21736, -313, 11191, -7981]
        --[0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0]
        (b"0000000000000000", b"0000000000000000", b"1001", b"0000", b"1111111111111111", b"00101010"),
        (b"0111111111111111", b"0000000000000000", b"1001", b"0000", b"0111111111111110", b"01010010"),
        (b"1000000000000000", b"0000000000000000", b"1001", b"0000", b"1011111111111111", b"10101010"),
        (b"0000000000000001", b"0000000000000000", b"1001", b"0000", b"0000000000000000", b"01100001"),
        (b"1101000100101100", b"0000000000000000", b"1001", b"0000", b"1101000100101011", b"00101010"),
        (b"1010100011101001", b"0000000000000000", b"1001", b"0000", b"1010100011101000", b"00101010"),
        (b"0101100100011110", b"0000000000000000", b"1001", b"0000", b"0101100100011101", b"01010010"),
        (b"1011011100111001", b"0000000000000000", b"1001", b"0000", b"1011011100111000", b"00101010"),
        (b"0111001010100110", b"0000000000000000", b"1001", b"0000", b"0111001010100101", b"01010010"),
        (b"0011101101000001", b"0000000000000000", b"1001", b"0000", b"0011101101000000", b"01010010"),
        (b"0000110100010010", b"0000000000000000", b"1001", b"0000", b"0000110100010001", b"01010010"),
        (b"1010101100011000", b"0000000000000000", b"1001", b"0000", b"1010101100010111", b"00101010"),
        (b"1111111011000111", b"0000000000000000", b"1001", b"0000", b"1111111011000110", b"00101010"),
        (b"0010101110110111", b"0000000000000000", b"1001", b"0000", b"0010101110110110", b"01010010"),
        (b"1110000011010011", b"0000000000000000", b"1001", b"0000", b"1110000011010010", b"00101010"),
        --A+B
        --[0, 32767, -32768, 1, 17050, -20330, 9253, -16612, 25346, -5742, -18759, 9089, -12291, -19773, 22974]
        --[18564, -12055, 30087, -4013, 12554, 15826, 27893, 11116, -32173, -6421, 24996, -31521, 23465, 9236, 21082]
        (b"0000000000000000", b"0100100010000100", b"1010", b"0000", b"0100100010000100", b"01010010"),
        (b"0111111111111111", b"1101000011101001", b"1010", b"0000", b"0101000011101000", b"01010010"),
        (b"1000000000000000", b"0111010110000111", b"1010", b"0000", b"1111010110000111", b"00101010"),
        (b"0000000000000001", b"1111000001010011", b"1010", b"0000", b"1111000001010100", b"00101010"),
        (b"0100001010011010", b"0011000100001010", b"1010", b"0000", b"0111001110100100", b"01010010"),
        (b"1011000010010110", b"0011110111010010", b"1010", b"0000", b"1110111001101000", b"00101010"),
        (b"0010010000100101", b"0110110011110101", b"1010", b"0000", b"1001000100011010", b"11010010"),
        (b"1011111100011100", b"0010101101101100", b"1010", b"0000", b"1110101010001000", b"00101010"),
        (b"0110001100000010", b"1000001001010011", b"1010", b"0000", b"1110010101010101", b"00101010"),
        (b"1110100110010010", b"1110011011101011", b"1010", b"0000", b"1101000001111101", b"00101010"),
        (b"1011011010111001", b"0110000110100100", b"1010", b"0000", b"0001100001011101", b"01010010"),
        (b"0010001110000001", b"1000010011011111", b"1010", b"0000", b"1010100001100000", b"00101010"),
        (b"1100111111111101", b"0101101110101001", b"1010", b"0000", b"0010101110100110", b"01010010"),
        (b"1011001011000011", b"0010010000010100", b"1010", b"0000", b"1101011011010111", b"00101010"),
        (b"0101100110111110", b"0101001001011010", b"1010", b"0000", b"1010110000011000", b"11010010"),
        --A-B
        --[0, 32767, -32768, 1, -20369, 8553, -21567, -32569, -87, 1745, -993, -8601, -14518, 21746, 22955]
        --[-14786, 8574, -13442, 10025, -7402, 5964, 28503, 27491, 15579, -2388, -30507, 9767, -3909, -18063, -28511]
        (b"0000000000000000", b"1100011000111110", b"1011", b"0000", b"0011100111000010", b"01010010"),
        (b"0111111111111111", b"0010000101111110", b"1011", b"0000", b"0101111010000001", b"01010010"),
        (b"1000000000000000", b"1100101101111110", b"1011", b"0000", b"1011010010000010", b"00101010"),
        (b"0000000000000001", b"0010011100101001", b"1011", b"0000", b"1101100011011000", b"00101010"),
        (b"1011000001101111", b"1110001100010110", b"1011", b"0000", b"1100110101011001", b"00101010"),
        (b"0010000101101001", b"0001011101001100", b"1011", b"0000", b"0000101000011101", b"01010010"),
        (b"1010101111000001", b"0110111101010111", b"1011", b"0000", b"1001111000110101", b"10101010"),
        (b"1000000011000111", b"0110101101100011", b"1011", b"0000", b"1000101010110010", b"10101010"),
        (b"1111111110101001", b"0011110011011011", b"1011", b"0000", b"1100001011001110", b"00101010"),
        (b"0000011011010001", b"1111011010101100", b"1011", b"0000", b"0001000000100101", b"01010010"),
        (b"1111110000011111", b"1000100011010101", b"1011", b"0000", b"0111001101001010", b"01010010"),
        (b"1101111001100111", b"0010011000100111", b"1011", b"0000", b"1011100001000000", b"00101010"),
        (b"1100011101001010", b"1111000010111011", b"1011", b"0000", b"1101011010001111", b"00101010"),
        (b"0101010011110010", b"1011100101110001", b"1011", b"0000", b"1001101110000001", b"11010010"),
        (b"0101100110101011", b"1001000010100001", b"1011", b"0000", b"1100100100001010", b"11010010"),
            --A<<SH
            --[1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1]
            --[0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0]
            (b"0000000000000001", b"0000000000000000", x"C", x"0", b"0000000000000001", b"01010110"),
            (b"0000000000000001", b"0000000000000000", x"C", x"1", b"0000000000000010", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"2", b"0000000000000100", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"3", b"0000000000001000", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"4", b"0000000000010000", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"5", b"0000000000100000", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"6", b"0000000001000000", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"7", b"0000000010000000", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"9", b"0000000100000000", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"A", b"0000010000000000", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"B", b"0000100000000000", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"C", b"0001000000000000", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"D", b"0010000000000000", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"E", b"0100000000000000", b"01010010"),
            (b"0000000000000001", b"0000000000000000", x"C", x"F", b"1000000000000000", b"00101010"),
            --A>>SH
            --[-32768, -32768, -32768, -32768, -32768, -32768, -32768, -32768, -32768, -32768, -32768, -32768, -32768, -32768, -32768, -32768]
            --[0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0]
            (b"1000000000000000", b"0000000000000000", x"D", x"0", b"1000000000000000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"1", b"1100000000000000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"2", b"1110000000000000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"3", b"1111000000000000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"4", b"1111100000000000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"5", b"1111110000000000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"6", b"1111111000000000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"7", b"1111111100000000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"8", b"1111111110000000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"9", b"1111111111000000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"A", b"1111111111100000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"B", b"1111111111110000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"C", b"1111111111111000", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"D", b"1111111111111100", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"E", b"1111111111111110", b"00101010"),
            (b"1000000000000000", b"0000000000000000", x"D", x"F", b"1111111111111111", b"00101010")
        );
begin

UUT : entity work.param_ALU
        generic map ( data_size => data_size)
        port map ( A => A, -- configure ports
                   B => B,
                   opcode => opcode,
                   SH => SH,
                   Output => Output,
                   flags => flags);
tb: process 
begin
    wait for 100ns;
    for i in test_vectors'range loop -- loop test vectors
        A <= test_vectors(i).A_TV; -- assign vector values
        B <= test_vectors(i).B_TV;
        opcode <= test_vectors(i).opcode_TV;
        SH <= test_vectors(i).SH_TV;
        Output <= test_vectors(i).Output_TV;
        flags <= test_vectors(i).flags_TV;
        wait for 20ns; -- allow propergation
        -- assert correct operation
        assert ((Output = test_vectors(i).Output_TV)
            and (flags = test_vectors(i).flags_TV))
        report -- if output doesn't match expected output
            "Test sequence " &
             integer'image(i+1) &
             " failed : " &
             " A is "&
             integer'image(to_integer(unsigned(A))) &
             " B is "&
             integer'image(to_integer(unsigned(B))) &
             ", opcode "&
             integer'image(to_integer(unsigned(opcode)))&
             ", ALU_output : "&
              integer'image(to_integer(unsigned(Output))) &
             ", expected : "&
              integer'image(to_integer(unsigned(test_vectors(i).Output_TV)))&
              ", ALU_flags : ZERO FLAG = "&
              std_logic'image(flags(0))&
              ", ZERO FLAG exp. = "&
              std_logic'image(test_vectors(i).flags_TV(0))&
              ", NON ZERO FLAG = "&
              std_logic'image(flags(1))&
              ", NON ZERO FLAG exp. = "&
              std_logic'image(test_vectors(i).flags_TV(1))&
              ", UNITY FLAG = "&
              std_logic'image(flags(2))&
              ", UNITY FLAG exp. = "&
              std_logic'image(test_vectors(i).flags_TV(2))&
              ", NEGATIVE FLAG = "&
              std_logic'image(flags(3))&
              ", NEGATIVE FLAG exp. = "&
              std_logic'image(test_vectors(i).flags_TV(3))&
              ", POSITIVE FLAG = "&
              std_logic'image(flags(4))&
              ", POSITIVE FLAG exp. = "&
              std_logic'image(test_vectors(i).flags_TV(4))&
              ", NON-POSITIVE FLAG = "&
              std_logic'image(flags(5))&
              ", NON-POSITIVE FLAG exp. = "&
              std_logic'image(test_vectors(i).flags_TV(5))&
              ", NON-NEGATIVE FLAG = "&
              std_logic'image(flags(6))&
              ", NON-NEGATIVE FLAG exp. = "&
              std_logic'image(test_vectors(i).flags_TV(6))&
              ", OVERFLOW FLAG = "&
              std_logic'image(flags(7))&
              ", OVERFLOW FLAG exp. = "&
              std_logic'image(test_vectors(i).flags_TV(7))
        severity note;
        end loop;
    wait;
end process;
end Behavioral;
